CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 140 1 200 9
0 71 1920 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
25 C:\CircuitMaker 6\BOM.DAT
0 7
0 71 1920 1040
143654930 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 201 559 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
2 +V
167 214 507 0 1 3
0 2
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
9 2-In AND~
219 381 414 0 3 22
0 9 5 11
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U4A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1132506026
65 0 0 0 4 1 4 0
1 U
3618 0 0
0
0
8 2-In OR~
219 400 356 0 3 22
0 11 10 8
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U3B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 -1300278184
65 0 0 0 4 2 3 0
1 U
6153 0 0
0
0
8 2-In OR~
219 271 425 0 3 22
0 4 13 12
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U3A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -1216392099
65 0 0 0 4 1 3 0
1 U
5394 0 0
0
0
7 Pulser~
4 540 524 0 10 12
0 15 16 14 17 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7734 0 0
0
0
14 Logic Display~
6 712 173 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 579 173 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 445 173 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 302 173 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
5 4027~
219 709 315 0 7 32
0 18 4 14 5 3 10 6
0
0 0 4720 90
4 4027
7 -60 35 -52
3 U2B
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 512 2 2 2 0
1 U
9325 0 0
0
0
5 4027~
219 578 314 0 7 32
0 3 6 14 7 19 4 5
0
0 0 4720 90
4 4027
7 -60 35 -52
3 U2A
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 512 2 1 2 0
1 U
8903 0 0
0
0
5 4027~
219 444 313 0 7 32
0 20 4 14 8 3 21 13
0
0 0 4720 90
4 4027
7 -60 35 -52
3 U1B
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 512 2 2 1 0
1 U
3834 0 0
0
0
5 4027~
219 295 311 0 7 32
0 22 12 14 2 3 7 9
0
0 0 4720 90
4 4027
7 -60 35 -52
3 U1A
33 -52 54 -44
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 975089484
65 0 0 512 2 1 1 0
1 U
3363 0 0
0
0
26
4 1 2 0 0 4224 0 14 2 0 0 3
306 312
306 516
214 516
5 0 3 0 0 8320 0 14 0 0 5 3
330 288
331 288
331 559
5 0 3 0 0 0 0 11 0 0 4 4
744 292
760 292
760 559
496 559
1 0 3 0 0 0 0 12 0 0 5 4
550 291
496 291
496 559
484 559
5 1 3 0 0 128 0 13 1 0 0 4
479 290
484 290
484 559
213 559
2 0 4 0 0 8192 0 11 0 0 18 3
702 316
702 320
638 320
0 4 5 0 0 8320 0 0 11 12 0 6
565 259
565 250
752 250
752 327
720 327
720 316
0 2 6 0 0 12416 0 0 12 26 0 5
702 258
748 258
748 323
571 323
571 315
4 6 7 0 0 8320 0 12 14 0 0 6
589 315
589 319
335 319
335 250
306 250
306 258
2 0 4 0 0 8192 0 13 0 0 18 3
437 314
437 331
638 331
4 3 8 0 0 8320 0 13 4 0 0 4
455 314
455 325
403 325
403 326
0 2 5 0 0 0 0 0 3 25 0 4
568 259
545 259
545 435
389 435
0 1 9 0 0 8320 0 0 3 23 0 4
288 255
357 255
357 435
371 435
6 2 10 0 0 12416 0 11 4 0 0 4
720 262
769 262
769 372
412 372
1 3 11 0 0 8320 0 4 3 0 0 4
394 372
394 383
380 383
380 390
2 3 12 0 0 4224 0 14 5 0 0 4
288 312
288 394
274 394
274 395
0 2 13 0 0 12416 0 0 5 24 0 4
437 253
506 253
506 441
283 441
6 1 4 0 0 12416 0 12 5 0 0 5
589 261
638 261
638 453
265 453
265 441
3 0 14 0 0 4096 0 13 0 0 22 2
446 314
446 469
3 0 14 0 0 0 0 12 0 0 22 2
580 315
580 469
3 0 14 0 0 0 0 11 0 0 22 2
711 316
711 469
3 3 14 0 0 8320 0 14 6 0 0 5
297 312
297 469
711 469
711 515
564 515
7 1 9 0 0 0 0 14 10 0 0 4
288 264
288 199
302 199
302 191
7 1 13 0 0 0 0 13 9 0 0 4
437 266
437 192
445 192
445 191
7 1 5 0 0 0 0 12 8 0 0 5
571 267
568 267
568 192
579 192
579 191
7 1 6 0 0 0 0 11 7 0 0 3
702 268
702 191
712 191
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
537 232 561 256
547 240 563 256
2 Q2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
671 222 695 246
681 230 697 246
2 Q3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
407 230 431 254
417 238 433 254
2 Q1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
253 242 277 266
263 250 279 266
2 QO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
182 566 262 590
192 574 264 590
9 Reiniciar
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
